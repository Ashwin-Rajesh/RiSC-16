/*
MIT License

Copyright (c) 2022 Ashwin Rajesh

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.
*/

`ifndef DESIGN_SV
`define DESIGN_SV

`include "core.v"

module toplevel (
  input clk,                  // Global clock
  output[15:0] pc
);

  localparam p_INST_NUM = 1024;
  localparam p_CODE_FILE = "code.data";
  
  reg[15:0] memory[p_INST_NUM];

  initial begin
    $readmemb(p_CODE_FILE, memory);
  end

  core #(.p_DATA_MEM_SIZE(1024)) processor_core (
      .clk(clk),
      .rst(0),
      .instruction(memory[pc]),
      .pc(pc)
  );
  
endmodule

`endif
